library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ff is
    	Port (
       		clk : in std_logic := '0';      
        	we  : in std_logic := '0';        
        	input   : in std_logic :='0'; 
        	output   : out std_logic := '0'
    	);
end ff;


architecture Behavioral of ff is
    	signal reg : std_logic := '0';
begin
    	process(clk)
    	begin
        	if rising_edge(clk) then
            		if we = '1' then
                		reg <= input;
            		end if;
        	end if;
    	end process;
    	output <= reg;
end Behavioral;
